-- megafunction wizard: %ALTSQRT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsqrt 

-- ============================================================
-- File Name: SqrRt32ClkEn.vhd
-- Megafunction Name(s):
-- 			altsqrt
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 5.1 Build 213 01/19/2006 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2006 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SqrRt32ClkEn IS
	PORT
	(
		clk		: IN STD_LOGIC ;
		ena		: IN STD_LOGIC ;
		radical		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		q		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		remainder		: OUT STD_LOGIC_VECTOR (16 DOWNTO 0)
	);
END SqrRt32ClkEn;


ARCHITECTURE SYN OF sqrrt32clken IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (16 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (15 DOWNTO 0);



	COMPONENT altsqrt
	GENERIC (
		pipeline		: NATURAL;
		q_port_width		: NATURAL;
		r_port_width		: NATURAL;
		width		: NATURAL;
		lpm_type		: STRING
	);
	PORT (
			remainder	: OUT STD_LOGIC_VECTOR (16 DOWNTO 0);
			radical	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ena	: IN STD_LOGIC ;
			q	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			clk	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	remainder    <= sub_wire0(16 DOWNTO 0);
	q    <= sub_wire1(15 DOWNTO 0);

	altsqrt_component : altsqrt
	GENERIC MAP (
		pipeline => 1,
		q_port_width => 16,
		r_port_width => 17,
		width => 32,
		lpm_type => "altsqrt"
	)
	PORT MAP (
		radical => radical,
		ena => ena,
		clk => clk,
		remainder => sub_wire0,
		q => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "1"
-- Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "16"
-- Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "17"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "32"
-- Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL clk
-- Retrieval info: USED_PORT: ena 0 0 0 0 INPUT NODEFVAL ena
-- Retrieval info: USED_PORT: q 0 0 16 0 OUTPUT NODEFVAL q[15..0]
-- Retrieval info: USED_PORT: radical 0 0 32 0 INPUT NODEFVAL radical[31..0]
-- Retrieval info: USED_PORT: remainder 0 0 17 0 OUTPUT NODEFVAL remainder[16..0]
-- Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
-- Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
-- Retrieval info: CONNECT: @radical 0 0 32 0 radical 0 0 32 0
-- Retrieval info: CONNECT: q 0 0 16 0 @q 0 0 16 0
-- Retrieval info: CONNECT: remainder 0 0 17 0 @remainder 0 0 17 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL SqrRt32ClkEn.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL SqrRt32ClkEn.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL SqrRt32ClkEn.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL SqrRt32ClkEn.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL SqrRt32ClkEn_inst.vhd FALSE
