/*=================================================================*\
Filename				:	dev_led.v
Author				:	Wisely
Description			:	
Revision	History	:	2017-04-07
							V1.0
Company				:
Email					:
Copyright(c) ,DreamFly Technology Inc,All right reserved
\*=================================================================*/
module dev_led(
	led
);

//============================================================
//Post in/out
//============================================================
output led;

//============================================================
//Assignment
//============================================================

assign led = 0;







endmodule
